module p1();


endmodule
