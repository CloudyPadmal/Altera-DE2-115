module Digitizer3(lineIns, LEDs);
	
	// Inputs and outputs
	input [7:0] lineIns;
	output [20:0] LEDs;
	
	reg [3:0] bcd0In;
	reg [3:0] bcd1In;
	reg [3:0] bcd2In;
	
	// Create two BCDs
	BCD bcd0(.lineIn(bcd0In), .lineOut(LEDs[6:0]));
	BCD bcd1(.lineIn(bcd1In), .lineOut(LEDs[13:7]));
	BCD bcd2(.lineIn(bcd2In), .lineOut(LEDs[20:14]));
	
	always @ *
		case (lineIns)
			8'b00000000 : begin bcd0In = 4'b0000; bcd1In = 4'b0000; bcd2In = 4'b0000; end // 00
			8'b00000001 : begin bcd0In = 4'b0001; bcd1In = 4'b0000; bcd2In = 4'b0000; end // 01
			8'b00000010 : begin bcd0In = 4'b0010; bcd1In = 4'b0000; bcd2In = 4'b0000; end // 02
			8'b00000011 : begin bcd0In = 4'b0011; bcd1In = 4'b0000; bcd2In = 4'b0000; end // 03
			8'b00000100 : begin bcd0In = 4'b0100; bcd1In = 4'b0000; bcd2In = 4'b0000; end // 04
			8'b00000101 : begin bcd0In = 4'b0101; bcd1In = 4'b0000; bcd2In = 4'b0000; end // 05
			8'b00000110 : begin bcd0In = 4'b0110; bcd1In = 4'b0000; bcd2In = 4'b0000; end // 06
			8'b00000111 : begin bcd0In = 4'b0111; bcd1In = 4'b0000; bcd2In = 4'b0000; end // 07
			8'b00001000 : begin bcd0In = 4'b1000; bcd1In = 4'b0000; bcd2In = 4'b0000; end // 08
			8'b00001001 : begin bcd0In = 4'b1000; bcd1In = 4'b0000; bcd2In = 4'b0000; end // 09
			8'b00001010 : begin bcd0In = 4'b0000; bcd1In = 4'b0001; bcd2In = 4'b0000; end // 10
			8'b00001011 : begin bcd0In = 4'b0001; bcd1In = 4'b0001; bcd2In = 4'b0000; end // 11
			8'b00001100 : begin bcd0In = 4'b0010; bcd1In = 4'b0001; bcd2In = 4'b0000; end // 12
			8'b00001101 : begin bcd0In = 4'b0011; bcd1In = 4'b0001; bcd2In = 4'b0000; end // 13
			8'b00001110 : begin bcd0In = 4'b0100; bcd1In = 4'b0001; bcd2In = 4'b0000; end // 14
			8'b00001111 : begin bcd0In = 4'b0101; bcd1In = 4'b0001; bcd2In = 4'b0000; end // 15
			8'b00010000 : begin bcd0In = 4'b0110; bcd1In = 4'b0001; bcd2In = 4'b0000; end // 16
			8'b00010001 : begin bcd0In = 4'b0111; bcd1In = 4'b0001; bcd2In = 4'b0000; end // 17
			8'b00010010 : begin bcd0In = 4'b1000; bcd1In = 4'b0001; bcd2In = 4'b0000; end // 18
			8'b00010011 : begin bcd0In = 4'b1001; bcd1In = 4'b0001; bcd2In = 4'b0000; end // 19
			8'b00010100 : begin bcd0In = 4'b0000; bcd1In = 4'b0010; bcd2In = 4'b0000; end // 20
			8'b00010101 : begin bcd0In = 4'b0001; bcd1In = 4'b0010; bcd2In = 4'b0000; end // 21
			8'b00010110 : begin bcd0In = 4'b0010; bcd1In = 4'b0010; bcd2In = 4'b0000; end // 22
			8'b00010111 : begin bcd0In = 4'b0011; bcd1In = 4'b0010; bcd2In = 4'b0000; end // 23
			8'b00011000 : begin bcd0In = 4'b0100; bcd1In = 4'b0010; bcd2In = 4'b0000; end // 24
			8'b00011001 : begin bcd0In = 4'b0101; bcd1In = 4'b0010; bcd2In = 4'b0000; end // 25
			8'b00011010 : begin bcd0In = 4'b0110; bcd1In = 4'b0010; bcd2In = 4'b0000; end // 26
			8'b00011011 : begin bcd0In = 4'b0111; bcd1In = 4'b0010; bcd2In = 4'b0000; end // 27
			8'b00011100 : begin bcd0In = 4'b1000; bcd1In = 4'b0010; bcd2In = 4'b0000; end // 28
			8'b00011101 : begin bcd0In = 4'b1001; bcd1In = 4'b0010; bcd2In = 4'b0000; end // 29
			8'b00011110 : begin bcd0In = 4'b0000; bcd1In = 4'b0011; bcd2In = 4'b0000; end // 30
			8'b00011111 : begin bcd0In = 4'b0001; bcd1In = 4'b0011; bcd2In = 4'b0000; end // 31
			8'b00100000 : begin bcd0In = 4'b0010; bcd1In = 4'b0011; bcd2In = 4'b0000; end // 32
			8'b00100001 : begin bcd0In = 4'b0011; bcd1In = 4'b0011; bcd2In = 4'b0000; end // 33
			8'b00100010 : begin bcd0In = 4'b0100; bcd1In = 4'b0011; bcd2In = 4'b0000; end // 34
			8'b00100011 : begin bcd0In = 4'b0101; bcd1In = 4'b0011; bcd2In = 4'b0000; end // 35
			8'b00100100 : begin bcd0In = 4'b0110; bcd1In = 4'b0011; bcd2In = 4'b0000; end // 36
			8'b00100101 : begin bcd0In = 4'b0111; bcd1In = 4'b0011; bcd2In = 4'b0000; end // 37
			8'b00100110 : begin bcd0In = 4'b1000; bcd1In = 4'b0011; bcd2In = 4'b0000; end // 38
			8'b00100111 : begin bcd0In = 4'b1001; bcd1In = 4'b0011; bcd2In = 4'b0000; end // 39
			8'b00101000 : begin bcd0In = 4'b0000; bcd1In = 4'b0100; bcd2In = 4'b0000; end // 40
			8'b00101001 : begin bcd0In = 4'b0001; bcd1In = 4'b0100; bcd2In = 4'b0000; end // 41
			8'b00101010 : begin bcd0In = 4'b0010; bcd1In = 4'b0100; bcd2In = 4'b0000; end // 42
			8'b00101011 : begin bcd0In = 4'b0011; bcd1In = 4'b0100; bcd2In = 4'b0000; end // 43
			8'b00101100 : begin bcd0In = 4'b0100; bcd1In = 4'b0100; bcd2In = 4'b0000; end // 44
			8'b00101101 : begin bcd0In = 4'b0101; bcd1In = 4'b0100; bcd2In = 4'b0000; end // 45
			8'b00101110 : begin bcd0In = 4'b0110; bcd1In = 4'b0100; bcd2In = 4'b0000; end // 46
			8'b00101111 : begin bcd0In = 4'b0111; bcd1In = 4'b0100; bcd2In = 4'b0000; end // 47
			8'b00110000 : begin bcd0In = 4'b1000; bcd1In = 4'b0100; bcd2In = 4'b0000; end // 48
			8'b00110001 : begin bcd0In = 4'b1001; bcd1In = 4'b0100; bcd2In = 4'b0000; end // 49
			8'b00110010 : begin bcd0In = 4'b0000; bcd1In = 4'b0101; bcd2In = 4'b0000; end // 50
			8'b00110011 : begin bcd0In = 4'b0001; bcd1In = 4'b0101; bcd2In = 4'b0000; end // 51
			8'b00110100 : begin bcd0In = 4'b0010; bcd1In = 4'b0101; bcd2In = 4'b0000; end // 52
			8'b00110101 : begin bcd0In = 4'b0011; bcd1In = 4'b0101; bcd2In = 4'b0000; end // 53
			8'b00110110 : begin bcd0In = 4'b0100; bcd1In = 4'b0101; bcd2In = 4'b0000; end // 54
			8'b00110111 : begin bcd0In = 4'b0101; bcd1In = 4'b0101; bcd2In = 4'b0000; end // 55
			8'b00111000 : begin bcd0In = 4'b0110; bcd1In = 4'b0101; bcd2In = 4'b0000; end // 56
			8'b00111001 : begin bcd0In = 4'b0111; bcd1In = 4'b0101; bcd2In = 4'b0000; end // 57
			8'b00111010 : begin bcd0In = 4'b1000; bcd1In = 4'b0101; bcd2In = 4'b0000; end // 58
			8'b00111011 : begin bcd0In = 4'b1001; bcd1In = 4'b0101; bcd2In = 4'b0000; end // 59
			8'b00111100 : begin bcd0In = 4'b0000; bcd1In = 4'b0110; bcd2In = 4'b0000; end // 60
			8'b00111101 : begin bcd0In = 4'b0001; bcd1In = 4'b0110; bcd2In = 4'b0000; end // 61
			8'b00111110 : begin bcd0In = 4'b0010; bcd1In = 4'b0110; bcd2In = 4'b0000; end // 62
			8'b00111111 : begin bcd0In = 4'b0011; bcd1In = 4'b0110; bcd2In = 4'b0000; end // 63
			8'b01000000 : begin bcd0In = 4'b0100; bcd1In = 4'b0110; bcd2In = 4'b0000; end // 64
			8'b01000001 : begin bcd0In = 4'b0101; bcd1In = 4'b0110; bcd2In = 4'b0000; end // 65
			8'b01000010 : begin bcd0In = 4'b0110; bcd1In = 4'b0110; bcd2In = 4'b0000; end // 66
			8'b01000011 : begin bcd0In = 4'b0111; bcd1In = 4'b0110; bcd2In = 4'b0000; end // 67
			8'b01000100 : begin bcd0In = 4'b1000; bcd1In = 4'b0110; bcd2In = 4'b0000; end // 68
			8'b01000101 : begin bcd0In = 4'b1001; bcd1In = 4'b0110; bcd2In = 4'b0000; end // 69
			8'b01000110 : begin bcd0In = 4'b0000; bcd1In = 4'b0111; bcd2In = 4'b0000; end // 70
			8'b01000111 : begin bcd0In = 4'b0001; bcd1In = 4'b0111; bcd2In = 4'b0000; end // 71
			8'b01001000 : begin bcd0In = 4'b0010; bcd1In = 4'b0111; bcd2In = 4'b0000; end // 72
			8'b01001001 : begin bcd0In = 4'b0011; bcd1In = 4'b0111; bcd2In = 4'b0000; end // 73
			8'b01001010 : begin bcd0In = 4'b0100; bcd1In = 4'b0111; bcd2In = 4'b0000; end // 74
			8'b01001011 : begin bcd0In = 4'b0101; bcd1In = 4'b0111; bcd2In = 4'b0000; end // 75
			8'b01001100 : begin bcd0In = 4'b0110; bcd1In = 4'b0111; bcd2In = 4'b0000; end // 76
			8'b01001101 : begin bcd0In = 4'b0111; bcd1In = 4'b0111; bcd2In = 4'b0000; end // 77
			8'b01001110 : begin bcd0In = 4'b1000; bcd1In = 4'b0111; bcd2In = 4'b0000; end // 78
			8'b01001111 : begin bcd0In = 4'b1001; bcd1In = 4'b0111; bcd2In = 4'b0000; end // 79
			8'b01010000 : begin bcd0In = 4'b0000; bcd1In = 4'b1000; bcd2In = 4'b0000; end // 80
			8'b01010001 : begin bcd0In = 4'b0001; bcd1In = 4'b1000; bcd2In = 4'b0000; end // 81
			8'b01010010 : begin bcd0In = 4'b0010; bcd1In = 4'b1000; bcd2In = 4'b0000; end // 82
			8'b01010011 : begin bcd0In = 4'b0011; bcd1In = 4'b1000; bcd2In = 4'b0000; end // 83
			8'b01010100 : begin bcd0In = 4'b0100; bcd1In = 4'b1000; bcd2In = 4'b0000; end // 84
			8'b01010101 : begin bcd0In = 4'b0101; bcd1In = 4'b1000; bcd2In = 4'b0000; end // 85
			8'b01010110 : begin bcd0In = 4'b0110; bcd1In = 4'b1000; bcd2In = 4'b0000; end // 86
			8'b01010111 : begin bcd0In = 4'b0111; bcd1In = 4'b1000; bcd2In = 4'b0000; end // 87
			8'b01011000 : begin bcd0In = 4'b1000; bcd1In = 4'b1000; bcd2In = 4'b0000; end // 88
			8'b01011001 : begin bcd0In = 4'b1001; bcd1In = 4'b1000; bcd2In = 4'b0000; end // 89
			8'b01011010 : begin bcd0In = 4'b0000; bcd1In = 4'b1001; bcd2In = 4'b0000; end // 90
			8'b01011011 : begin bcd0In = 4'b0001; bcd1In = 4'b1001; bcd2In = 4'b0000; end // 91
			8'b01011100 : begin bcd0In = 4'b0010; bcd1In = 4'b1001; bcd2In = 4'b0000; end // 92
			8'b01011101 : begin bcd0In = 4'b0011; bcd1In = 4'b1001; bcd2In = 4'b0000; end // 93
			8'b01011110 : begin bcd0In = 4'b0100; bcd1In = 4'b1001; bcd2In = 4'b0000; end // 94
			8'b01011111 : begin bcd0In = 4'b0101; bcd1In = 4'b1001; bcd2In = 4'b0000; end // 95
			8'b01100000 : begin bcd0In = 4'b0110; bcd1In = 4'b1001; bcd2In = 4'b0000; end // 96
			8'b01100001 : begin bcd0In = 4'b0111; bcd1In = 4'b1001; bcd2In = 4'b0000; end // 97
			8'b01100010 : begin bcd0In = 4'b1000; bcd1In = 4'b1001; bcd2In = 4'b0000; end // 98
			8'b01100011 : begin bcd0In = 4'b1001; bcd1In = 4'b1001; bcd2In = 4'b0000; end // 99		
			8'b01100100 : begin bcd0In = 4'b0000; bcd1In = 4'b0000; bcd2In = 4'b0001; end // 100
			8'b01100101 : begin bcd0In = 4'b0001; bcd1In = 4'b0000; bcd2In = 4'b0001; end // 101
			8'b01100110 : begin bcd0In = 4'b0010; bcd1In = 4'b0000; bcd2In = 4'b0001; end // 102
			8'b01100111 : begin bcd0In = 4'b0011; bcd1In = 4'b0000; bcd2In = 4'b0001; end // 103
			8'b01101000 : begin bcd0In = 4'b0100; bcd1In = 4'b0000; bcd2In = 4'b0001; end // 104
			8'b01101001 : begin bcd0In = 4'b0101; bcd1In = 4'b0000; bcd2In = 4'b0001; end // 105
			8'b01101010 : begin bcd0In = 4'b0110; bcd1In = 4'b0000; bcd2In = 4'b0001; end // 106
			8'b01101011 : begin bcd0In = 4'b0111; bcd1In = 4'b0000; bcd2In = 4'b0001; end // 107
			8'b01101100 : begin bcd0In = 4'b1000; bcd1In = 4'b0000; bcd2In = 4'b0001; end // 108
			8'b01101101 : begin bcd0In = 4'b1001; bcd1In = 4'b0000; bcd2In = 4'b0001; end // 109
			8'b01101110 : begin bcd0In = 4'b0000; bcd1In = 4'b0001; bcd2In = 4'b0001; end // 110
			8'b01101111 : begin bcd0In = 4'b0001; bcd1In = 4'b0001; bcd2In = 4'b0001; end // 111
			8'b01110000 : begin bcd0In = 4'b0010; bcd1In = 4'b0001; bcd2In = 4'b0001; end // 112
			8'b01110001 : begin bcd0In = 4'b0011; bcd1In = 4'b0001; bcd2In = 4'b0001; end // 113
			8'b01110010 : begin bcd0In = 4'b0100; bcd1In = 4'b0001; bcd2In = 4'b0001; end // 114
			8'b01110011 : begin bcd0In = 4'b0101; bcd1In = 4'b0001; bcd2In = 4'b0001; end // 115
			8'b01110100 : begin bcd0In = 4'b0110; bcd1In = 4'b0001; bcd2In = 4'b0001; end // 116
			8'b01110101 : begin bcd0In = 4'b0111; bcd1In = 4'b0001; bcd2In = 4'b0001; end // 117
			8'b01110110 : begin bcd0In = 4'b1000; bcd1In = 4'b0001; bcd2In = 4'b0001; end // 118
			8'b01110111 : begin bcd0In = 4'b1001; bcd1In = 4'b0001; bcd2In = 4'b0001; end // 119
			8'b01111000 : begin bcd0In = 4'b0000; bcd1In = 4'b0010; bcd2In = 4'b0001; end // 120
			8'b01111001 : begin bcd0In = 4'b0001; bcd1In = 4'b0010; bcd2In = 4'b0001; end // 121
			8'b01111010 : begin bcd0In = 4'b0010; bcd1In = 4'b0010; bcd2In = 4'b0001; end // 122
			8'b01111011 : begin bcd0In = 4'b0011; bcd1In = 4'b0010; bcd2In = 4'b0001; end // 123
			8'b01111100 : begin bcd0In = 4'b0100; bcd1In = 4'b0010; bcd2In = 4'b0001; end // 124
			8'b01111101 : begin bcd0In = 4'b0101; bcd1In = 4'b0010; bcd2In = 4'b0001; end // 125
			8'b01111110 : begin bcd0In = 4'b0110; bcd1In = 4'b0010; bcd2In = 4'b0001; end // 126
			8'b01111111 : begin bcd0In = 4'b0111; bcd1In = 4'b0010; bcd2In = 4'b0001; end // 127
			8'b10000000 : begin bcd0In = 4'b1000; bcd1In = 4'b0010; bcd2In = 4'b0001; end // 128
			8'b10000001 : begin bcd0In = 4'b1001; bcd1In = 4'b0010; bcd2In = 4'b0001; end // 129
			8'b10000010 : begin bcd0In = 4'b0000; bcd1In = 4'b0011; bcd2In = 4'b0001; end // 130
			8'b10000011 : begin bcd0In = 4'b0001; bcd1In = 4'b0011; bcd2In = 4'b0001; end // 131
			8'b10000100 : begin bcd0In = 4'b0010; bcd1In = 4'b0011; bcd2In = 4'b0001; end // 132
			8'b10000101 : begin bcd0In = 4'b0011; bcd1In = 4'b0011; bcd2In = 4'b0001; end // 133
			8'b10000110 : begin bcd0In = 4'b0100; bcd1In = 4'b0011; bcd2In = 4'b0001; end // 134
			8'b10000111 : begin bcd0In = 4'b0101; bcd1In = 4'b0011; bcd2In = 4'b0001; end // 135
			8'b10001000 : begin bcd0In = 4'b0110; bcd1In = 4'b0011; bcd2In = 4'b0001; end // 136
			8'b10001001 : begin bcd0In = 4'b0111; bcd1In = 4'b0011; bcd2In = 4'b0001; end // 137
			8'b10001010 : begin bcd0In = 4'b1000; bcd1In = 4'b0011; bcd2In = 4'b0001; end // 138
			8'b10001011 : begin bcd0In = 4'b1001; bcd1In = 4'b0011; bcd2In = 4'b0001; end // 139
			8'b10001100 : begin bcd0In = 4'b0000; bcd1In = 4'b0100; bcd2In = 4'b0001; end // 140
			8'b10001101 : begin bcd0In = 4'b0001; bcd1In = 4'b0100; bcd2In = 4'b0001; end // 141
			8'b10001110 : begin bcd0In = 4'b0010; bcd1In = 4'b0100; bcd2In = 4'b0001; end // 142
			8'b10001111 : begin bcd0In = 4'b0011; bcd1In = 4'b0100; bcd2In = 4'b0001; end // 143
			8'b10010000 : begin bcd0In = 4'b0100; bcd1In = 4'b0100; bcd2In = 4'b0001; end // 144
			8'b10010001 : begin bcd0In = 4'b0101; bcd1In = 4'b0100; bcd2In = 4'b0001; end // 145
			8'b10010010 : begin bcd0In = 4'b0110; bcd1In = 4'b0100; bcd2In = 4'b0001; end // 146
			8'b10010011 : begin bcd0In = 4'b0111; bcd1In = 4'b0100; bcd2In = 4'b0001; end // 147
			8'b10010100 : begin bcd0In = 4'b1000; bcd1In = 4'b0100; bcd2In = 4'b0001; end // 148
			8'b10010101 : begin bcd0In = 4'b1001; bcd1In = 4'b0100; bcd2In = 4'b0001; end // 149
			8'b10010110 : begin bcd0In = 4'b0000; bcd1In = 4'b0101; bcd2In = 4'b0001; end // 150
			8'b10010111 : begin bcd0In = 4'b0001; bcd1In = 4'b0101; bcd2In = 4'b0001; end // 151
			8'b10011000 : begin bcd0In = 4'b0010; bcd1In = 4'b0101; bcd2In = 4'b0001; end // 152
			8'b10011001 : begin bcd0In = 4'b0011; bcd1In = 4'b0101; bcd2In = 4'b0001; end // 153
			8'b10011010 : begin bcd0In = 4'b0100; bcd1In = 4'b0101; bcd2In = 4'b0001; end // 154
			8'b10011011 : begin bcd0In = 4'b0101; bcd1In = 4'b0101; bcd2In = 4'b0001; end // 155
			8'b10011100 : begin bcd0In = 4'b0110; bcd1In = 4'b0101; bcd2In = 4'b0001; end // 156
			8'b10011101 : begin bcd0In = 4'b0111; bcd1In = 4'b0101; bcd2In = 4'b0001; end // 157
			8'b10011110 : begin bcd0In = 4'b1000; bcd1In = 4'b0101; bcd2In = 4'b0001; end // 158
			8'b10011111 : begin bcd0In = 4'b1001; bcd1In = 4'b0101; bcd2In = 4'b0001; end // 159
			8'b10100000 : begin bcd0In = 4'b0000; bcd1In = 4'b0110; bcd2In = 4'b0001; end // 160
			8'b10100001 : begin bcd0In = 4'b0001; bcd1In = 4'b0110; bcd2In = 4'b0001; end // 161
			8'b10100010 : begin bcd0In = 4'b0010; bcd1In = 4'b0110; bcd2In = 4'b0001; end // 162
			8'b10100011 : begin bcd0In = 4'b0011; bcd1In = 4'b0110; bcd2In = 4'b0001; end // 163
			8'b10100100 : begin bcd0In = 4'b0100; bcd1In = 4'b0110; bcd2In = 4'b0001; end // 164
			8'b10100101 : begin bcd0In = 4'b0101; bcd1In = 4'b0110; bcd2In = 4'b0001; end // 165
			8'b10100110 : begin bcd0In = 4'b0110; bcd1In = 4'b0110; bcd2In = 4'b0001; end // 166
			8'b10100111 : begin bcd0In = 4'b0111; bcd1In = 4'b0110; bcd2In = 4'b0001; end // 167
			8'b10101000 : begin bcd0In = 4'b1000; bcd1In = 4'b0110; bcd2In = 4'b0001; end // 168
			8'b10101001 : begin bcd0In = 4'b1001; bcd1In = 4'b0110; bcd2In = 4'b0001; end // 169
			8'b10101010 : begin bcd0In = 4'b0000; bcd1In = 4'b0111; bcd2In = 4'b0001; end // 170
			8'b10101011 : begin bcd0In = 4'b0001; bcd1In = 4'b0111; bcd2In = 4'b0001; end // 171
			8'b10101100 : begin bcd0In = 4'b0010; bcd1In = 4'b0111; bcd2In = 4'b0001; end // 172
			8'b10101101 : begin bcd0In = 4'b0011; bcd1In = 4'b0111; bcd2In = 4'b0001; end // 173
			8'b10101110 : begin bcd0In = 4'b0100; bcd1In = 4'b0111; bcd2In = 4'b0001; end // 174
			8'b10101111 : begin bcd0In = 4'b0101; bcd1In = 4'b0111; bcd2In = 4'b0001; end // 175
			8'b10110000 : begin bcd0In = 4'b0110; bcd1In = 4'b0111; bcd2In = 4'b0001; end // 176
			8'b10110001 : begin bcd0In = 4'b0111; bcd1In = 4'b0111; bcd2In = 4'b0001; end // 177
			8'b10110010 : begin bcd0In = 4'b1000; bcd1In = 4'b0111; bcd2In = 4'b0001; end // 178
			8'b10110011 : begin bcd0In = 4'b1001; bcd1In = 4'b0111; bcd2In = 4'b0001; end // 179
			8'b10110100 : begin bcd0In = 4'b0000; bcd1In = 4'b1000; bcd2In = 4'b0001; end // 180
			8'b10110101 : begin bcd0In = 4'b0001; bcd1In = 4'b1000; bcd2In = 4'b0001; end // 181
			8'b10110110 : begin bcd0In = 4'b0010; bcd1In = 4'b1000; bcd2In = 4'b0001; end // 182
			8'b10110111 : begin bcd0In = 4'b0011; bcd1In = 4'b1000; bcd2In = 4'b0001; end // 183
			8'b10111000 : begin bcd0In = 4'b0100; bcd1In = 4'b1000; bcd2In = 4'b0001; end // 184
			8'b10111001 : begin bcd0In = 4'b0101; bcd1In = 4'b1000; bcd2In = 4'b0001; end // 185
			8'b10111010 : begin bcd0In = 4'b0110; bcd1In = 4'b1000; bcd2In = 4'b0001; end // 186
			8'b10111011 : begin bcd0In = 4'b0111; bcd1In = 4'b1000; bcd2In = 4'b0001; end // 187
			8'b10111100 : begin bcd0In = 4'b1000; bcd1In = 4'b1000; bcd2In = 4'b0001; end // 188
			8'b10111101 : begin bcd0In = 4'b1001; bcd1In = 4'b1000; bcd2In = 4'b0001; end // 189
			8'b10111110 : begin bcd0In = 4'b0000; bcd1In = 4'b1001; bcd2In = 4'b0001; end // 190
			8'b10111111 : begin bcd0In = 4'b0001; bcd1In = 4'b1001; bcd2In = 4'b0001; end // 191
			8'b11000000 : begin bcd0In = 4'b0010; bcd1In = 4'b1001; bcd2In = 4'b0001; end // 192
			8'b11000001 : begin bcd0In = 4'b0011; bcd1In = 4'b1001; bcd2In = 4'b0001; end // 193
			8'b11000010 : begin bcd0In = 4'b0100; bcd1In = 4'b1001; bcd2In = 4'b0001; end // 194
			8'b11000011 : begin bcd0In = 4'b0101; bcd1In = 4'b1001; bcd2In = 4'b0001; end // 195
			8'b11000100 : begin bcd0In = 4'b0110; bcd1In = 4'b1001; bcd2In = 4'b0001; end // 196
			8'b11000101 : begin bcd0In = 4'b0111; bcd1In = 4'b1001; bcd2In = 4'b0001; end // 197
			8'b11000110 : begin bcd0In = 4'b1000; bcd1In = 4'b1001; bcd2In = 4'b0001; end // 198
			8'b11000111 : begin bcd0In = 4'b1001; bcd1In = 4'b1001; bcd2In = 4'b0001; end // 199
			default 		: begin bcd0In = 4'b0000; bcd1In = 4'b0000; bcd2In = 4'b0000; end
		endcase
endmodule